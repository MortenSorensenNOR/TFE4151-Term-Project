*.PARAM ln_or=0.2u   ! Length of NMOS transistors
*.PARAM wn_or=0.25u    ! Width  of NMOS transistors
*.PARAM lp_or=0.2u   ! Length of PMOS transistors
*.PARAM wp_or=1u    ! Width  of PMOS transistors

.PARAM ln_or=ln   ! Length of NMOS transistors
.PARAM wn_or=wn    ! Width  of NMOS transistors
.PARAM lp_or=lp   ! Length of PMOS transistors
.PARAM wp_or=wp    ! Width  of PMOS transistors

.subckt OR_GATE A B Y VDD VSS

* drain gate source bulk  <-- port order both n and p
* Pull-up network (PMOS transistors in series)
xmn1 T    A VDD VDD pmos1v l=lp_or w=wp_or      ! PMOS controlled by input A
xmn2 Yinv B T   T   pmos1v l=lp_or w=wp_or      ! PMOS controlled by input B (in series with xmn1)

* Pull-down network (NMOS transistors in series)
xmn3 Yinv A VSS VSS nmos1v l=ln_or w=wn_or   ! NMOS controlled by input A
xmn4 Yinv B VSS VSS nmos1v l=ln_or w=wn_or   ! NMOS controlled by input B (in paralell with xmn3)

* output inverter
xmn5 Y Yinv VDD VDD pmos1v l=lp_or w=wp_or   ! PMOS controlled by input Yinverted
xmn6 Y Yinv VSS VSS nmos1v l=ln_or w=wn_or   ! NMOS controlled by input Yinverted


.ends